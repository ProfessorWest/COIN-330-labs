module testlab02;

wire out;
wire nout;
reg in1;
lab02 testing(in1, out, nout);

initial begin

	in1 = 1'b0;
	#1 $display("in1=%b, out=%b, nout=%b", in1, out, nout);

	end
endmodule
